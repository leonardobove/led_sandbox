// led_sandbox_sopc.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module led_sandbox_sopc (
		inout  wire        accelerometer_spi_I2C_SDAT,      //  accelerometer_spi.I2C_SDAT
		output wire        accelerometer_spi_I2C_SCLK,      //                   .I2C_SCLK
		output wire        accelerometer_spi_G_SENSOR_CS_N, //                   .G_SENSOR_CS_N
		input  wire        accelerometer_spi_G_SENSOR_INT,  //                   .G_SENSOR_INT
		input  wire        clk_clk,                         //                clk.clk
		output wire        clk_sdram_clk,                   //          clk_sdram.clk
		output wire        led_matrix_clock_clk,            //   led_matrix_clock.clk
		output wire        led_matrix_control_row_sel_a,    // led_matrix_control.row_sel_a
		output wire        led_matrix_control_row_sel_b,    //                   .row_sel_b
		output wire        led_matrix_control_blue_1,       //                   .blue_1
		output wire        led_matrix_control_blue_2,       //                   .blue_2
		output wire        led_matrix_control_row_sel_c,    //                   .row_sel_c
		output wire        led_matrix_control_row_sel_d,    //                   .row_sel_d
		output wire        led_matrix_control_green_1,      //                   .green_1
		output wire        led_matrix_control_green_2,      //                   .green_2
		output wire        led_matrix_control_latch,        //                   .latch
		output wire        led_matrix_control_output_en,    //                   .output_en
		output wire        led_matrix_control_red_1,        //                   .red_1
		output wire        led_matrix_control_red_2,        //                   .red_2
		input  wire        reset_reset_n,                   //              reset.reset_n
		output wire [12:0] sdram_wire_addr,                 //         sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                   //                   .ba
		output wire        sdram_wire_cas_n,                //                   .cas_n
		output wire        sdram_wire_cke,                  //                   .cke
		output wire        sdram_wire_cs_n,                 //                   .cs_n
		inout  wire [15:0] sdram_wire_dq,                   //                   .dq
		output wire [1:0]  sdram_wire_dqm,                  //                   .dqm
		output wire        sdram_wire_ras_n,                //                   .ras_n
		output wire        sdram_wire_we_n                  //                   .we_n
	);

	wire         video_dma_controller_0_avalon_pixel_source_valid;                                      // video_dma_controller_0:stream_valid -> led_matrix_driver_0:valid
	wire  [15:0] video_dma_controller_0_avalon_pixel_source_data;                                       // video_dma_controller_0:stream_data -> led_matrix_driver_0:data
	wire         video_dma_controller_0_avalon_pixel_source_ready;                                      // led_matrix_driver_0:ready -> video_dma_controller_0:stream_ready
	wire         video_dma_controller_0_avalon_pixel_source_startofpacket;                              // video_dma_controller_0:stream_startofpacket -> led_matrix_driver_0:startofpacket
	wire         video_dma_controller_0_avalon_pixel_source_endofpacket;                                // video_dma_controller_0:stream_endofpacket -> led_matrix_driver_0:endofpacket
	wire         altpll_0_c0_clk;                                                                       // altpll_0:c0 -> [cpu:clk, irq_mapper:clk, irq_synchronizer:sender_clk, jtag_uart:clk, mm_interconnect_0:altpll_0_c0_clk, rst_controller_002:clk, sdram:clk, system_id:clock, systick_timer:clk]
	wire         altpll_0_c2_clk;                                                                       // altpll_0:c2 -> [accelerometer_spi_0:clk, irq_synchronizer:receiver_clk, mm_interconnect_0:altpll_0_c2_clk, rst_controller:clk]
	wire         altpll_0_c3_clk;                                                                       // altpll_0:c3 -> [led_matrix_driver_0:clock, mm_interconnect_0:altpll_0_c3_clk, rst_controller_003:clk, video_dma_controller_0:clk]
	wire         video_dma_controller_0_avalon_dma_master_waitrequest;                                  // mm_interconnect_0:video_dma_controller_0_avalon_dma_master_waitrequest -> video_dma_controller_0:master_waitrequest
	wire  [15:0] video_dma_controller_0_avalon_dma_master_readdata;                                     // mm_interconnect_0:video_dma_controller_0_avalon_dma_master_readdata -> video_dma_controller_0:master_readdata
	wire  [31:0] video_dma_controller_0_avalon_dma_master_address;                                      // video_dma_controller_0:master_address -> mm_interconnect_0:video_dma_controller_0_avalon_dma_master_address
	wire         video_dma_controller_0_avalon_dma_master_read;                                         // video_dma_controller_0:master_read -> mm_interconnect_0:video_dma_controller_0_avalon_dma_master_read
	wire         video_dma_controller_0_avalon_dma_master_readdatavalid;                                // mm_interconnect_0:video_dma_controller_0_avalon_dma_master_readdatavalid -> video_dma_controller_0:master_readdatavalid
	wire         video_dma_controller_0_avalon_dma_master_lock;                                         // video_dma_controller_0:master_arbiterlock -> mm_interconnect_0:video_dma_controller_0_avalon_dma_master_lock
	wire  [31:0] cpu_data_master_readdata;                                                              // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                                           // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                                           // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [27:0] cpu_data_master_address;                                                               // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                                            // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                                                  // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_write;                                                                 // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                                             // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                                                       // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                                                    // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [27:0] cpu_instruction_master_address;                                                        // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                                           // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         mm_interconnect_0_sdram_s1_chipselect;                                                 // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                                                   // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                                                // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                                                    // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                                       // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                                                 // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                                              // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                                      // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                                                  // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;                                        // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;                                     // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;                                     // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;                                         // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                                            // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;                                      // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;                                           // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;                                       // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire   [7:0] mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_readdata;    // accelerometer_spi_0:readdata -> mm_interconnect_0:accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_readdata
	wire         mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_waitrequest; // accelerometer_spi_0:waitrequest -> mm_interconnect_0:accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_waitrequest
	wire   [0:0] mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_address;     // mm_interconnect_0:accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_address -> accelerometer_spi_0:address
	wire         mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_read;        // mm_interconnect_0:accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_read -> accelerometer_spi_0:read
	wire   [0:0] mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_byteenable;  // mm_interconnect_0:accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_byteenable -> accelerometer_spi_0:byteenable
	wire         mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_write;       // mm_interconnect_0:accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_write -> accelerometer_spi_0:write
	wire   [7:0] mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_writedata;   // mm_interconnect_0:accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_writedata -> accelerometer_spi_0:writedata
	wire  [31:0] mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_readdata;            // video_dma_controller_0:slave_readdata -> mm_interconnect_0:video_dma_controller_0_avalon_dma_control_slave_readdata
	wire   [1:0] mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_address;             // mm_interconnect_0:video_dma_controller_0_avalon_dma_control_slave_address -> video_dma_controller_0:slave_address
	wire         mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_read;                // mm_interconnect_0:video_dma_controller_0_avalon_dma_control_slave_read -> video_dma_controller_0:slave_read
	wire   [3:0] mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_byteenable;          // mm_interconnect_0:video_dma_controller_0_avalon_dma_control_slave_byteenable -> video_dma_controller_0:slave_byteenable
	wire         mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_write;               // mm_interconnect_0:video_dma_controller_0_avalon_dma_control_slave_write -> video_dma_controller_0:slave_write
	wire  [31:0] mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_writedata;           // mm_interconnect_0:video_dma_controller_0_avalon_dma_control_slave_writedata -> video_dma_controller_0:slave_writedata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;                              // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                                // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;                             // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                                 // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                                    // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                                   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_led_matrix_driver_0_avalon_slave_0_readdata;                         // led_matrix_driver_0:readdata -> mm_interconnect_0:led_matrix_driver_0_avalon_slave_0_readdata
	wire   [0:0] mm_interconnect_0_led_matrix_driver_0_avalon_slave_0_address;                          // mm_interconnect_0:led_matrix_driver_0_avalon_slave_0_address -> led_matrix_driver_0:address
	wire         mm_interconnect_0_led_matrix_driver_0_avalon_slave_0_read;                             // mm_interconnect_0:led_matrix_driver_0_avalon_slave_0_read -> led_matrix_driver_0:read
	wire         mm_interconnect_0_led_matrix_driver_0_avalon_slave_0_write;                            // mm_interconnect_0:led_matrix_driver_0_avalon_slave_0_write -> led_matrix_driver_0:write
	wire  [31:0] mm_interconnect_0_led_matrix_driver_0_avalon_slave_0_writedata;                        // mm_interconnect_0:led_matrix_driver_0_avalon_slave_0_writedata -> led_matrix_driver_0:writedata
	wire  [31:0] mm_interconnect_0_system_id_control_slave_readdata;                                    // system_id:readdata -> mm_interconnect_0:system_id_control_slave_readdata
	wire   [0:0] mm_interconnect_0_system_id_control_slave_address;                                     // mm_interconnect_0:system_id_control_slave_address -> system_id:address
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_readdata;                                         // altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_0_pll_slave_address;                                          // mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	wire         mm_interconnect_0_altpll_0_pll_slave_read;                                             // mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	wire         mm_interconnect_0_altpll_0_pll_slave_write;                                            // mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_writedata;                                        // mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	wire         mm_interconnect_0_systick_timer_s1_chipselect;                                         // mm_interconnect_0:systick_timer_s1_chipselect -> systick_timer:chipselect
	wire  [15:0] mm_interconnect_0_systick_timer_s1_readdata;                                           // systick_timer:readdata -> mm_interconnect_0:systick_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_systick_timer_s1_address;                                            // mm_interconnect_0:systick_timer_s1_address -> systick_timer:address
	wire         mm_interconnect_0_systick_timer_s1_write;                                              // mm_interconnect_0:systick_timer_s1_write -> systick_timer:write_n
	wire  [15:0] mm_interconnect_0_systick_timer_s1_writedata;                                          // mm_interconnect_0:systick_timer_s1_writedata -> systick_timer:writedata
	wire         irq_mapper_receiver1_irq;                                                              // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                              // systick_timer:irq -> irq_mapper:receiver2_irq
	wire  [31:0] cpu_irq_irq;                                                                           // irq_mapper:sender_irq -> cpu:irq
	wire         irq_mapper_receiver0_irq;                                                              // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                                         // accelerometer_spi_0:irq -> irq_synchronizer:receiver_irq
	wire         rst_controller_reset_out_reset;                                                        // rst_controller:reset_out -> [accelerometer_spi_0:reset, irq_synchronizer:receiver_reset, mm_interconnect_0:accelerometer_spi_0_reset_reset_bridge_in_reset_reset]
	wire         cpu_debug_reset_request_reset;                                                         // cpu:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in1]
	wire         rst_controller_001_reset_out_reset;                                                    // rst_controller_001:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_002_reset_out_reset;                                                    // rst_controller_002:reset_out -> [cpu:reset_n, irq_mapper:reset, irq_synchronizer:sender_reset, jtag_uart:rst_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, sdram:reset_n, system_id:reset_n, systick_timer:reset_n]
	wire         rst_controller_002_reset_out_reset_req;                                                // rst_controller_002:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_003_reset_out_reset;                                                    // rst_controller_003:reset_out -> [led_matrix_driver_0:areset_n, mm_interconnect_0:video_dma_controller_0_reset_reset_bridge_in_reset_reset, video_dma_controller_0:reset]

	led_sandbox_sopc_accelerometer_spi_0 accelerometer_spi_0 (
		.clk           (altpll_0_c2_clk),                                                                       //                                 clk.clk
		.reset         (rst_controller_reset_out_reset),                                                        //                               reset.reset
		.address       (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_address),     // avalon_accelerometer_spi_mode_slave.address
		.byteenable    (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_byteenable),  //                                    .byteenable
		.read          (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_read),        //                                    .read
		.write         (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_write),       //                                    .write
		.writedata     (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_writedata),   //                                    .writedata
		.readdata      (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_readdata),    //                                    .readdata
		.waitrequest   (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_waitrequest), //                                    .waitrequest
		.irq           (irq_synchronizer_receiver_irq),                                                         //                           interrupt.irq
		.I2C_SDAT      (accelerometer_spi_I2C_SDAT),                                                            //                  external_interface.export
		.I2C_SCLK      (accelerometer_spi_I2C_SCLK),                                                            //                                    .export
		.G_SENSOR_CS_N (accelerometer_spi_G_SENSOR_CS_N),                                                       //                                    .export
		.G_SENSOR_INT  (accelerometer_spi_G_SENSOR_INT)                                                         //                                    .export
	);

	led_sandbox_sopc_altpll_0 altpll_0 (
		.clk                (clk_clk),                                        //       inclk_interface.clk
		.reset              (rst_controller_001_reset_out_reset),             // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_0_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_0_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_0_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_0_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_0_pll_slave_writedata), //                      .writedata
		.c0                 (altpll_0_c0_clk),                                //                    c0.clk
		.c1                 (clk_sdram_clk),                                  //                    c1.clk
		.c2                 (altpll_0_c2_clk),                                //                    c2.clk
		.c3                 (altpll_0_c3_clk),                                //                    c3.clk
		.scandone           (),                                               //           (terminated)
		.scandataout        (),                                               //           (terminated)
		.c4                 (),                                               //           (terminated)
		.areset             (1'b0),                                           //           (terminated)
		.locked             (),                                               //           (terminated)
		.phasedone          (),                                               //           (terminated)
		.phasecounterselect (3'b000),                                         //           (terminated)
		.phaseupdown        (1'b0),                                           //           (terminated)
		.phasestep          (1'b0),                                           //           (terminated)
		.scanclk            (1'b0),                                           //           (terminated)
		.scanclkena         (1'b0),                                           //           (terminated)
		.scandata           (1'b0),                                           //           (terminated)
		.configupdate       (1'b0)                                            //           (terminated)
	);

	led_sandbox_sopc_cpu cpu (
		.clk                                 (altpll_0_c0_clk),                                   //                       clk.clk
		.reset_n                             (~rst_controller_002_reset_out_reset),               //                     reset.reset_n
		.reset_req                           (rst_controller_002_reset_out_reset_req),            //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	led_sandbox_sopc_jtag_uart jtag_uart (
		.clk            (altpll_0_c0_clk),                                           //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	led_matrix_driver #(
		.ENABLE_DEFAULT (1),
		.RESET_DEFAULT  (0),
		.MAT_WIDTH      (64),
		.MAT_HEIGHT     (32)
	) led_matrix_driver_0 (
		.address       (mm_interconnect_0_led_matrix_driver_0_avalon_slave_0_address),   //        avalon_slave_0.address
		.write         (mm_interconnect_0_led_matrix_driver_0_avalon_slave_0_write),     //                      .write
		.writedata     (mm_interconnect_0_led_matrix_driver_0_avalon_slave_0_writedata), //                      .writedata
		.readdata      (mm_interconnect_0_led_matrix_driver_0_avalon_slave_0_readdata),  //                      .readdata
		.read          (mm_interconnect_0_led_matrix_driver_0_avalon_slave_0_read),      //                      .read
		.ready         (video_dma_controller_0_avalon_pixel_source_ready),               // avalon_streaming_sink.ready
		.valid         (video_dma_controller_0_avalon_pixel_source_valid),               //                      .valid
		.data          (video_dma_controller_0_avalon_pixel_source_data),                //                      .data
		.startofpacket (video_dma_controller_0_avalon_pixel_source_startofpacket),       //                      .startofpacket
		.endofpacket   (video_dma_controller_0_avalon_pixel_source_endofpacket),         //                      .endofpacket
		.CLK           (led_matrix_clock_clk),                                           //             clock_out.clk
		.clock         (altpll_0_c3_clk),                                                //              clock_in.clk
		.areset_n      (~rst_controller_003_reset_out_reset),                            //                 reset.reset_n
		.A             (led_matrix_control_row_sel_a),                                   //           conduit_out.row_sel_a
		.B             (led_matrix_control_row_sel_b),                                   //                      .row_sel_b
		.B1            (led_matrix_control_blue_1),                                      //                      .blue_1
		.B2            (led_matrix_control_blue_2),                                      //                      .blue_2
		.C             (led_matrix_control_row_sel_c),                                   //                      .row_sel_c
		.D             (led_matrix_control_row_sel_d),                                   //                      .row_sel_d
		.G1            (led_matrix_control_green_1),                                     //                      .green_1
		.G2            (led_matrix_control_green_2),                                     //                      .green_2
		.LAT           (led_matrix_control_latch),                                       //                      .latch
		.OE_n          (led_matrix_control_output_en),                                   //                      .output_en
		.R1            (led_matrix_control_red_1),                                       //                      .red_1
		.R2            (led_matrix_control_red_2)                                        //                      .red_2
	);

	led_sandbox_sopc_sdram sdram (
		.clk            (altpll_0_c0_clk),                          //   clk.clk
		.reset_n        (~rst_controller_002_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	led_sandbox_sopc_system_id system_id (
		.clock    (altpll_0_c0_clk),                                    //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_system_id_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_system_id_control_slave_address)   //              .address
	);

	led_sandbox_sopc_systick_timer systick_timer (
		.clk        (altpll_0_c0_clk),                               //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),           // reset.reset_n
		.address    (mm_interconnect_0_systick_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_systick_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_systick_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_systick_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_systick_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                       //   irq.irq
	);

	led_sandbox_sopc_video_dma_controller_0 video_dma_controller_0 (
		.clk                  (altpll_0_c3_clk),                                                              //                      clk.clk
		.reset                (rst_controller_003_reset_out_reset),                                           //                    reset.reset
		.master_address       (video_dma_controller_0_avalon_dma_master_address),                             //        avalon_dma_master.address
		.master_waitrequest   (video_dma_controller_0_avalon_dma_master_waitrequest),                         //                         .waitrequest
		.master_arbiterlock   (video_dma_controller_0_avalon_dma_master_lock),                                //                         .lock
		.master_read          (video_dma_controller_0_avalon_dma_master_read),                                //                         .read
		.master_readdata      (video_dma_controller_0_avalon_dma_master_readdata),                            //                         .readdata
		.master_readdatavalid (video_dma_controller_0_avalon_dma_master_readdatavalid),                       //                         .readdatavalid
		.slave_address        (mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_address),    // avalon_dma_control_slave.address
		.slave_byteenable     (mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_byteenable), //                         .byteenable
		.slave_read           (mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_read),       //                         .read
		.slave_write          (mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_write),      //                         .write
		.slave_writedata      (mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_writedata),  //                         .writedata
		.slave_readdata       (mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_readdata),   //                         .readdata
		.stream_ready         (video_dma_controller_0_avalon_pixel_source_ready),                             //      avalon_pixel_source.ready
		.stream_data          (video_dma_controller_0_avalon_pixel_source_data),                              //                         .data
		.stream_startofpacket (video_dma_controller_0_avalon_pixel_source_startofpacket),                     //                         .startofpacket
		.stream_endofpacket   (video_dma_controller_0_avalon_pixel_source_endofpacket),                       //                         .endofpacket
		.stream_valid         (video_dma_controller_0_avalon_pixel_source_valid)                              //                         .valid
	);

	led_sandbox_sopc_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c0_clk                                                     (altpll_0_c0_clk),                                                                       //                                             altpll_0_c0.clk
		.altpll_0_c2_clk                                                     (altpll_0_c2_clk),                                                                       //                                             altpll_0_c2.clk
		.altpll_0_c3_clk                                                     (altpll_0_c3_clk),                                                                       //                                             altpll_0_c3.clk
		.clk_50_clk_clk                                                      (clk_clk),                                                                               //                                              clk_50_clk.clk
		.accelerometer_spi_0_reset_reset_bridge_in_reset_reset               (rst_controller_reset_out_reset),                                                        //         accelerometer_spi_0_reset_reset_bridge_in_reset.reset
		.altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset          (rst_controller_001_reset_out_reset),                                                    //    altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
		.cpu_reset_reset_bridge_in_reset_reset                               (rst_controller_002_reset_out_reset),                                                    //                         cpu_reset_reset_bridge_in_reset.reset
		.video_dma_controller_0_reset_reset_bridge_in_reset_reset            (rst_controller_003_reset_out_reset),                                                    //      video_dma_controller_0_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                                             (cpu_data_master_address),                                                               //                                         cpu_data_master.address
		.cpu_data_master_waitrequest                                         (cpu_data_master_waitrequest),                                                           //                                                        .waitrequest
		.cpu_data_master_byteenable                                          (cpu_data_master_byteenable),                                                            //                                                        .byteenable
		.cpu_data_master_read                                                (cpu_data_master_read),                                                                  //                                                        .read
		.cpu_data_master_readdata                                            (cpu_data_master_readdata),                                                              //                                                        .readdata
		.cpu_data_master_write                                               (cpu_data_master_write),                                                                 //                                                        .write
		.cpu_data_master_writedata                                           (cpu_data_master_writedata),                                                             //                                                        .writedata
		.cpu_data_master_debugaccess                                         (cpu_data_master_debugaccess),                                                           //                                                        .debugaccess
		.cpu_instruction_master_address                                      (cpu_instruction_master_address),                                                        //                                  cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                                  (cpu_instruction_master_waitrequest),                                                    //                                                        .waitrequest
		.cpu_instruction_master_read                                         (cpu_instruction_master_read),                                                           //                                                        .read
		.cpu_instruction_master_readdata                                     (cpu_instruction_master_readdata),                                                       //                                                        .readdata
		.video_dma_controller_0_avalon_dma_master_address                    (video_dma_controller_0_avalon_dma_master_address),                                      //                video_dma_controller_0_avalon_dma_master.address
		.video_dma_controller_0_avalon_dma_master_waitrequest                (video_dma_controller_0_avalon_dma_master_waitrequest),                                  //                                                        .waitrequest
		.video_dma_controller_0_avalon_dma_master_read                       (video_dma_controller_0_avalon_dma_master_read),                                         //                                                        .read
		.video_dma_controller_0_avalon_dma_master_readdata                   (video_dma_controller_0_avalon_dma_master_readdata),                                     //                                                        .readdata
		.video_dma_controller_0_avalon_dma_master_readdatavalid              (video_dma_controller_0_avalon_dma_master_readdatavalid),                                //                                                        .readdatavalid
		.video_dma_controller_0_avalon_dma_master_lock                       (video_dma_controller_0_avalon_dma_master_lock),                                         //                                                        .lock
		.accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_address     (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_address),     // accelerometer_spi_0_avalon_accelerometer_spi_mode_slave.address
		.accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_write       (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_write),       //                                                        .write
		.accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_read        (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_read),        //                                                        .read
		.accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_readdata    (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_readdata),    //                                                        .readdata
		.accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_writedata   (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_writedata),   //                                                        .writedata
		.accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_byteenable  (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_byteenable),  //                                                        .byteenable
		.accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_waitrequest (mm_interconnect_0_accelerometer_spi_0_avalon_accelerometer_spi_mode_slave_waitrequest), //                                                        .waitrequest
		.altpll_0_pll_slave_address                                          (mm_interconnect_0_altpll_0_pll_slave_address),                                          //                                      altpll_0_pll_slave.address
		.altpll_0_pll_slave_write                                            (mm_interconnect_0_altpll_0_pll_slave_write),                                            //                                                        .write
		.altpll_0_pll_slave_read                                             (mm_interconnect_0_altpll_0_pll_slave_read),                                             //                                                        .read
		.altpll_0_pll_slave_readdata                                         (mm_interconnect_0_altpll_0_pll_slave_readdata),                                         //                                                        .readdata
		.altpll_0_pll_slave_writedata                                        (mm_interconnect_0_altpll_0_pll_slave_writedata),                                        //                                                        .writedata
		.cpu_debug_mem_slave_address                                         (mm_interconnect_0_cpu_debug_mem_slave_address),                                         //                                     cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                                           (mm_interconnect_0_cpu_debug_mem_slave_write),                                           //                                                        .write
		.cpu_debug_mem_slave_read                                            (mm_interconnect_0_cpu_debug_mem_slave_read),                                            //                                                        .read
		.cpu_debug_mem_slave_readdata                                        (mm_interconnect_0_cpu_debug_mem_slave_readdata),                                        //                                                        .readdata
		.cpu_debug_mem_slave_writedata                                       (mm_interconnect_0_cpu_debug_mem_slave_writedata),                                       //                                                        .writedata
		.cpu_debug_mem_slave_byteenable                                      (mm_interconnect_0_cpu_debug_mem_slave_byteenable),                                      //                                                        .byteenable
		.cpu_debug_mem_slave_waitrequest                                     (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),                                     //                                                        .waitrequest
		.cpu_debug_mem_slave_debugaccess                                     (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),                                     //                                                        .debugaccess
		.jtag_uart_avalon_jtag_slave_address                                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),                                 //                             jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                                   //                                                        .write
		.jtag_uart_avalon_jtag_slave_read                                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                                    //                                                        .read
		.jtag_uart_avalon_jtag_slave_readdata                                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),                                //                                                        .readdata
		.jtag_uart_avalon_jtag_slave_writedata                               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),                               //                                                        .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),                             //                                                        .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),                              //                                                        .chipselect
		.led_matrix_driver_0_avalon_slave_0_address                          (mm_interconnect_0_led_matrix_driver_0_avalon_slave_0_address),                          //                      led_matrix_driver_0_avalon_slave_0.address
		.led_matrix_driver_0_avalon_slave_0_write                            (mm_interconnect_0_led_matrix_driver_0_avalon_slave_0_write),                            //                                                        .write
		.led_matrix_driver_0_avalon_slave_0_read                             (mm_interconnect_0_led_matrix_driver_0_avalon_slave_0_read),                             //                                                        .read
		.led_matrix_driver_0_avalon_slave_0_readdata                         (mm_interconnect_0_led_matrix_driver_0_avalon_slave_0_readdata),                         //                                                        .readdata
		.led_matrix_driver_0_avalon_slave_0_writedata                        (mm_interconnect_0_led_matrix_driver_0_avalon_slave_0_writedata),                        //                                                        .writedata
		.sdram_s1_address                                                    (mm_interconnect_0_sdram_s1_address),                                                    //                                                sdram_s1.address
		.sdram_s1_write                                                      (mm_interconnect_0_sdram_s1_write),                                                      //                                                        .write
		.sdram_s1_read                                                       (mm_interconnect_0_sdram_s1_read),                                                       //                                                        .read
		.sdram_s1_readdata                                                   (mm_interconnect_0_sdram_s1_readdata),                                                   //                                                        .readdata
		.sdram_s1_writedata                                                  (mm_interconnect_0_sdram_s1_writedata),                                                  //                                                        .writedata
		.sdram_s1_byteenable                                                 (mm_interconnect_0_sdram_s1_byteenable),                                                 //                                                        .byteenable
		.sdram_s1_readdatavalid                                              (mm_interconnect_0_sdram_s1_readdatavalid),                                              //                                                        .readdatavalid
		.sdram_s1_waitrequest                                                (mm_interconnect_0_sdram_s1_waitrequest),                                                //                                                        .waitrequest
		.sdram_s1_chipselect                                                 (mm_interconnect_0_sdram_s1_chipselect),                                                 //                                                        .chipselect
		.system_id_control_slave_address                                     (mm_interconnect_0_system_id_control_slave_address),                                     //                                 system_id_control_slave.address
		.system_id_control_slave_readdata                                    (mm_interconnect_0_system_id_control_slave_readdata),                                    //                                                        .readdata
		.systick_timer_s1_address                                            (mm_interconnect_0_systick_timer_s1_address),                                            //                                        systick_timer_s1.address
		.systick_timer_s1_write                                              (mm_interconnect_0_systick_timer_s1_write),                                              //                                                        .write
		.systick_timer_s1_readdata                                           (mm_interconnect_0_systick_timer_s1_readdata),                                           //                                                        .readdata
		.systick_timer_s1_writedata                                          (mm_interconnect_0_systick_timer_s1_writedata),                                          //                                                        .writedata
		.systick_timer_s1_chipselect                                         (mm_interconnect_0_systick_timer_s1_chipselect),                                         //                                                        .chipselect
		.video_dma_controller_0_avalon_dma_control_slave_address             (mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_address),             //         video_dma_controller_0_avalon_dma_control_slave.address
		.video_dma_controller_0_avalon_dma_control_slave_write               (mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_write),               //                                                        .write
		.video_dma_controller_0_avalon_dma_control_slave_read                (mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_read),                //                                                        .read
		.video_dma_controller_0_avalon_dma_control_slave_readdata            (mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_readdata),            //                                                        .readdata
		.video_dma_controller_0_avalon_dma_control_slave_writedata           (mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_writedata),           //                                                        .writedata
		.video_dma_controller_0_avalon_dma_control_slave_byteenable          (mm_interconnect_0_video_dma_controller_0_avalon_dma_control_slave_byteenable)           //                                                        .byteenable
	);

	led_sandbox_sopc_irq_mapper irq_mapper (
		.clk           (altpll_0_c0_clk),                    //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.sender_irq    (cpu_irq_irq)                         //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (altpll_0_c2_clk),                    //       receiver_clk.clk
		.sender_clk     (altpll_0_c0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),  // reset_in1.reset
		.clk            (altpll_0_c2_clk),                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),          // reset_in1.reset
		.clk            (altpll_0_c0_clk),                        //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (altpll_0_c3_clk),                    //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
